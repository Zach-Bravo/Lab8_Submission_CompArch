module ROM(addr, dout);

input [31:0] addr;
output reg [31:0] dout;

always@(addr) begin
	case(addr)
		32'd00: dout = 32'b0;
	   32'd04: dout = 32'b00000000100000000000011010010011; //4 addi x13,x0,8 fixed
		32'd08: dout = 32'b00000000110101110010000000100011; //8 sw x13, 0(x14)
																			  //     rs2,imm/rs2,rs1
		32'd12: dout = 32'b00000000110101110010100000000011; //12 lw x16,0(x14) check				  
		//00000000010000000000011010010011	
		/*32'd08: dout = 32'b0;	
      32'd12: dout = 32'b00000000110101110010000000100011; //8 sw x13, 0(x14)
		32'd16: dout = 32'b00000000000001110010100000000011; //12 lw x16,0(x14) check
		//32'd04: dout = 32'b101101110110010001100011; //8 lw x5,x0,9*/		
		//32'd04: dout = 32'b101101110110010001100011; //8 lw x5,x0,9*/
		/*32'd00: dout = 32'h00450693; //0 addi x5,x0,9
		32'd04: dout = 32'h00100713; //4
		32'd08: dout = 32'h00b76463; //8
		32'd12: dout = 32'h00008067; //c
		32'd16: dout = 32'h0006a803; //10
		32'd20: dout = 32'h00068613; //14
		32'd24: dout = 32'h00070793; //18
		32'd28: dout = 32'hffc62883; //1c
		32'd32: dout = 32'h01185a63; //20
		32'd36: dout = 32'h01162023; //24
		32'd40: dout = 32'hfff78793; //28
		32'd44: dout = 32'hffc60613; //2c
		32'd48: dout = 32'hfe0796e3; //30
		32'd52: dout = 32'h00279793; //34
		32'd56: dout = 32'h00f507b3; //38
		32'd60: dout = 32'h0107a023; //3c
		32'd64: dout = 32'h00170713; //40
		32'd68: dout = 32'h00468693; //44
		32'd72: dout = 32'hfc1ff06f; //48*/
	
		default: dout = 32'd0;

	endcase 
end

endmodule 